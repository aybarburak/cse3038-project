module control(in,regdest,alusrc,memtoreg,regwrite,memread,memwrite,branch,bmve,balne,jalpce,bleze,bneale,balrne,aluop4,aluop3,aluop1,aluop2,select_ori,instruct,ne);
input [5:0] in,instruct;
output regdest,alusrc,memtoreg,regwrite,memread,memwrite,branch,balne,jalpce,aluop1,aluop2,aluop3,aluop4,select_ori,bleze,bneale,balrne,bmve,ne;
wire rformat,lw,sw,beq,bmv,baln,jalpc,ori,blez,bneal,balrn,ne;
assign rformat=~|in;
assign lw=in[5]& (~in[4])&(~in[3])&(~in[2])&in[1]&in[0];
assign sw=in[5]& (~in[4])&in[3]&(~in[2])&in[1]&in[0];
assign beq=~in[5]& (~in[4])&(~in[3])&in[2]&(~in[1])&(~in[0]);
assign bmv=(~in[5])& in[4]&(~in[3])&in[2]&in[1]&(~in[0]);
assign baln=in[5]& (~in[4])&(~in[3])&(~in[2])&(~in[1])&(~in[0]);
assign jalpc=(~in[5])& in[4]&in[3]&in[2]&in[1]&in[0];
assign ori=(~in[5])& (~in[4])&in[3]&in[2]&(~in[1])&in[0];
assign blez=(~in[5])& (~in[4])&(~in[3])&in[2]&in[1]&(~in[0]);
assign bneal=in[5]& (~in[4])&in[3]&in[2]&(~in[1])&in[0];
assign balrn=(~instruct[5])& instruct[4]&instruct[3]&(~instruct[2])&(~instruct[1])&(~instruct[0]);
assign regdest=rformat|balrn;
assign alusrc=lw|sw|bmv|ori;
assign memtoreg=lw;
assign regwrite=rformat|lw|baln|jalpc|ori|(bneal&ne)|balrn;
assign memread=lw|bmv;
assign memwrite=sw;
assign branch=beq;
assign bmve=bmv;
assign balne=baln;
assign jalpce=jalpc;
assign bleze=blez;
assign bneale=bneal;
assign balrne=balrn;
assign aluop1=rformat;
assign aluop2=beq;
assign aluop3=bmv;
assign aluop4=ori;
assign select_ori=ori;
endmodule
